`default_nettype none

module sine_lut (
  input  wire [7:0] addr,        // phase input (0–255)
  output reg  [7:0] amplitude    // corresponding sine amplitude
);

  always @(*) begin
    case (addr)
      8'd0: amplitude = 8'd128;
      8'd1: amplitude = 8'd131;
      8'd2: amplitude = 8'd134;
      8'd3: amplitude = 8'd137;
      8'd4: amplitude = 8'd140;
      8'd5: amplitude = 8'd143;
      8'd6: amplitude = 8'd146;
      8'd7: amplitude = 8'd149;
      8'd8: amplitude = 8'd152;
      8'd9: amplitude = 8'd155;
      8'd10: amplitude = 8'd158;
      8'd11: amplitude = 8'd162;
      8'd12: amplitude = 8'd165;
      8'd13: amplitude = 8'd167;
      8'd14: amplitude = 8'd170;
      8'd15: amplitude = 8'd173;
      8'd16: amplitude = 8'd176;
      8'd17: amplitude = 8'd179;
      8'd18: amplitude = 8'd182;
      8'd19: amplitude = 8'd185;
      8'd20: amplitude = 8'd188;
      8'd21: amplitude = 8'd190;
      8'd22: amplitude = 8'd193;
      8'd23: amplitude = 8'd196;
      8'd24: amplitude = 8'd198;
      8'd25: amplitude = 8'd201;
      8'd26: amplitude = 8'd203;
      8'd27: amplitude = 8'd206;
      8'd28: amplitude = 8'd208;
      8'd29: amplitude = 8'd211;
      8'd30: amplitude = 8'd213;
      8'd31: amplitude = 8'd215;
      8'd32: amplitude = 8'd218;
      8'd33: amplitude = 8'd220;
      8'd34: amplitude = 8'd222;
      8'd35: amplitude = 8'd224;
      8'd36: amplitude = 8'd226;
      8'd37: amplitude = 8'd228;
      8'd38: amplitude = 8'd230;
      8'd39: amplitude = 8'd232;
      8'd40: amplitude = 8'd234;
      8'd41: amplitude = 8'd235;
      8'd42: amplitude = 8'd237;
      8'd43: amplitude = 8'd238;
      8'd44: amplitude = 8'd240;
      8'd45: amplitude = 8'd241;
      8'd46: amplitude = 8'd243;
      8'd47: amplitude = 8'd244;
      8'd48: amplitude = 8'd245;
      8'd49: amplitude = 8'd246;
      8'd50: amplitude = 8'd248;
      8'd51: amplitude = 8'd249;
      8'd52: amplitude = 8'd250;
      8'd53: amplitude = 8'd250;
      8'd54: amplitude = 8'd251;
      8'd55: amplitude = 8'd252;
      8'd56: amplitude = 8'd253;
      8'd57: amplitude = 8'd253;
      8'd58: amplitude = 8'd254;
      8'd59: amplitude = 8'd254;
      8'd60: amplitude = 8'd254;
      8'd61: amplitude = 8'd255;
      8'd62: amplitude = 8'd255;
      8'd63: amplitude = 8'd255;
      8'd64: amplitude = 8'd255;
      8'd65: amplitude = 8'd255;
      8'd66: amplitude = 8'd255;
      8'd67: amplitude = 8'd255;
      8'd68: amplitude = 8'd254;
      8'd69: amplitude = 8'd254;
      8'd70: amplitude = 8'd254;
      8'd71: amplitude = 8'd253;
      8'd72: amplitude = 8'd253;
      8'd73: amplitude = 8'd252;
      8'd74: amplitude = 8'd251;
      8'd75: amplitude = 8'd250;
      8'd76: amplitude = 8'd250;
      8'd77: amplitude = 8'd249;
      8'd78: amplitude = 8'd248;
      8'd79: amplitude = 8'd246;
      8'd80: amplitude = 8'd245;
      8'd81: amplitude = 8'd244;
      8'd82: amplitude = 8'd243;
      8'd83: amplitude = 8'd241;
      8'd84: amplitude = 8'd240;
      8'd85: amplitude = 8'd238;
      8'd86: amplitude = 8'd237;
      8'd87: amplitude = 8'd235;
      8'd88: amplitude = 8'd234;
      8'd89: amplitude = 8'd232;
      8'd90: amplitude = 8'd230;
      8'd91: amplitude = 8'd228;
      8'd92: amplitude = 8'd226;
      8'd93: amplitude = 8'd224;
      8'd94: amplitude = 8'd222;
      8'd95: amplitude = 8'd220;
      8'd96: amplitude = 8'd218;
      8'd97: amplitude = 8'd215;
      8'd98: amplitude = 8'd213;
      8'd99: amplitude = 8'd211;
      8'd100: amplitude = 8'd208;
      8'd101: amplitude = 8'd206;
      8'd102: amplitude = 8'd203;
      8'd103: amplitude = 8'd201;
      8'd104: amplitude = 8'd198;
      8'd105: amplitude = 8'd196;
      8'd106: amplitude = 8'd193;
      8'd107: amplitude = 8'd190;
      8'd108: amplitude = 8'd188;
      8'd109: amplitude = 8'd185;
      8'd110: amplitude = 8'd182;
      8'd111: amplitude = 8'd179;
      8'd112: amplitude = 8'd176;
      8'd113: amplitude = 8'd173;
      8'd114: amplitude = 8'd170;
      8'd115: amplitude = 8'd167;
      8'd116: amplitude = 8'd165;
      8'd117: amplitude = 8'd162;
      8'd118: amplitude = 8'd158;
      8'd119: amplitude = 8'd155;
      8'd120: amplitude = 8'd152;
      8'd121: amplitude = 8'd149;
      8'd122: amplitude = 8'd146;
      8'd123: amplitude = 8'd143;
      8'd124: amplitude = 8'd140;
      8'd125: amplitude = 8'd137;
      8'd126: amplitude = 8'd134;
      8'd127: amplitude = 8'd131;
      8'd128: amplitude = 8'd128;
      8'd129: amplitude = 8'd124;
      8'd130: amplitude = 8'd121;
      8'd131: amplitude = 8'd118;
      8'd132: amplitude = 8'd115;
      8'd133: amplitude = 8'd112;
      8'd134: amplitude = 8'd109;
      8'd135: amplitude = 8'd106;
      8'd136: amplitude = 8'd103;
      8'd137: amplitude = 8'd100;
      8'd138: amplitude = 8'd97;
      8'd139: amplitude = 8'd93;
      8'd140: amplitude = 8'd90;
      8'd141: amplitude = 8'd88;
      8'd142: amplitude = 8'd85;
      8'd143: amplitude = 8'd82;
      8'd144: amplitude = 8'd79;
      8'd145: amplitude = 8'd76;
      8'd146: amplitude = 8'd73;
      8'd147: amplitude = 8'd70;
      8'd148: amplitude = 8'd67;
      8'd149: amplitude = 8'd65;
      8'd150: amplitude = 8'd62;
      8'd151: amplitude = 8'd59;
      8'd152: amplitude = 8'd57;
      8'd153: amplitude = 8'd54;
      8'd154: amplitude = 8'd52;
      8'd155: amplitude = 8'd49;
      8'd156: amplitude = 8'd47;
      8'd157: amplitude = 8'd44;
      8'd158: amplitude = 8'd42;
      8'd159: amplitude = 8'd40;
      8'd160: amplitude = 8'd37;
      8'd161: amplitude = 8'd35;
      8'd162: amplitude = 8'd33;
      8'd163: amplitude = 8'd31;
      8'd164: amplitude = 8'd29;
      8'd165: amplitude = 8'd27;
      8'd166: amplitude = 8'd25;
      8'd167: amplitude = 8'd23;
      8'd168: amplitude = 8'd21;
      8'd169: amplitude = 8'd20;
      8'd170: amplitude = 8'd18;
      8'd171: amplitude = 8'd17;
      8'd172: amplitude = 8'd15;
      8'd173: amplitude = 8'd14;
      8'd174: amplitude = 8'd12;
      8'd175: amplitude = 8'd11;
      8'd176: amplitude = 8'd10;
      8'd177: amplitude = 8'd9;
      8'd178: amplitude = 8'd7;
      8'd179: amplitude = 8'd6;
      8'd180: amplitude = 8'd5;
      8'd181: amplitude = 8'd5;
      8'd182: amplitude = 8'd4;
      8'd183: amplitude = 8'd3;
      8'd184: amplitude = 8'd2;
      8'd185: amplitude = 8'd2;
      8'd186: amplitude = 8'd1;
      8'd187: amplitude = 8'd1;
      8'd188: amplitude = 8'd1;
      8'd189: amplitude = 8'd0;
      8'd190: amplitude = 8'd0;
      8'd191: amplitude = 8'd0;
      8'd192: amplitude = 8'd0;
      8'd193: amplitude = 8'd0;
      8'd194: amplitude = 8'd0;
      8'd195: amplitude = 8'd0;
      8'd196: amplitude = 8'd1;
      8'd197: amplitude = 8'd1;
      8'd198: amplitude = 8'd1;
      8'd199: amplitude = 8'd2;
      8'd200: amplitude = 8'd2;
      8'd201: amplitude = 8'd3;
      8'd202: amplitude = 8'd4;
      8'd203: amplitude = 8'd5;
      8'd204: amplitude = 8'd5;
      8'd205: amplitude = 8'd6;
      8'd206: amplitude = 8'd7;
      8'd207: amplitude = 8'd9;
      8'd208: amplitude = 8'd10;
      8'd209: amplitude = 8'd11;
      8'd210: amplitude = 8'd12;
      8'd211: amplitude = 8'd14;
      8'd212: amplitude = 8'd15;
      8'd213: amplitude = 8'd17;
      8'd214: amplitude = 8'd18;
      8'd215: amplitude = 8'd20;
      8'd216: amplitude = 8'd21;
      8'd217: amplitude = 8'd23;
      8'd218: amplitude = 8'd25;
      8'd219: amplitude = 8'd27;
      8'd220: amplitude = 8'd29;
      8'd221: amplitude = 8'd31;
      8'd222: amplitude = 8'd33;
      8'd223: amplitude = 8'd35;
      8'd224: amplitude = 8'd37;
      8'd225: amplitude = 8'd40;
      8'd226: amplitude = 8'd42;
      8'd227: amplitude = 8'd44;
      8'd228: amplitude = 8'd47;
      8'd229: amplitude = 8'd49;
      8'd230: amplitude = 8'd52;
      8'd231: amplitude = 8'd54;
      8'd232: amplitude = 8'd57;
      8'd233: amplitude = 8'd59;
      8'd234: amplitude = 8'd62;
      8'd235: amplitude = 8'd65;
      8'd236: amplitude = 8'd67;
      8'd237: amplitude = 8'd70;
      8'd238: amplitude = 8'd73;
      8'd239: amplitude = 8'd76;
      8'd240: amplitude = 8'd79;
      8'd241: amplitude = 8'd82;
      8'd242: amplitude = 8'd85;
      8'd243: amplitude = 8'd88;
      8'd244: amplitude = 8'd90;
      8'd245: amplitude = 8'd93;
      8'd246: amplitude = 8'd97;
      8'd247: amplitude = 8'd100;
      8'd248: amplitude = 8'd103;
      8'd249: amplitude = 8'd106;
      8'd250: amplitude = 8'd109;
      8'd251: amplitude = 8'd112;
      8'd252: amplitude = 8'd115;
      8'd253: amplitude = 8'd118;
      8'd254: amplitude = 8'd121;
      8'd255: amplitude = 8'd124;
      default: amplitude = 8'd128;
    endcase
  end

endmodule
